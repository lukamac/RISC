library ieee;
use ieee.std_logic_1164.all;

entity IF_stage is
	port(
		clk		: in std_logic;
		rst		: in std_logic
		
	);
	
end IF_stage;

architecture rtl of IF_stage is

begin


end rtl;

