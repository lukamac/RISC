use work.RISC_const_and_types.all;

package op_codes is
    constant ADD : op_t := "00000";
    constant SUB : op_t := "00001";
end package op_codes;
