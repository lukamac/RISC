library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.RISC_const_and_types.all;
use work.op_codes.all;


entity EX_stage is
    port
    (
        clk, rst    : in std_logic;

        -- Operation code
        ctrl_op     : in op_t;

        -- ALU input B signals
        b           : in word_t;
        pc_in       : in address_t;
        ctrl_alu_b  : in std_logic;

        -- ALU input C signals
        c, imm      : in word_t;
        ctrl_alu_c  : in std_logic;

        status           : out status_t;
        pc_out           : out address_t;
        alu_res, mdr_out : out word_t
    );
end entity EX_stage;


architecture rtl of EX_stage is

    component alu is
        port
        (
            op   : in op_t;
            b, c : in word_t;

            a    : out word_t
        );
    end component alu;

    signal ctrl_op_reg : op_t;
    signal imm_reg, b_reg, c_reg, pc_reg : word_t;
    signal alu_b, alu_c : word_t;

begin

    process (clk) is
    begin
        if (rising_edge(clk)) then
            if (rst = '1') then
                ctrl_op_reg <= (others => '0');
                imm_reg     <= (others => '0');
                b_reg       <= (others => '0');
                c_reg       <= (others => '0');
                pc_reg      <= (others => '0');
            else
                ctrl_op_reg <= ctrl_op;
                imm_reg     <= imm;
                b_reg       <= b;
                c_reg       <= c;
                pc_reg      <= pc;
            end if;
        end if;
    end process;

    alu_inst : component alu port map (op => ctrl_op_reg,
                                       b  => alu_b,
                                       c  => alu_c,
                                       a  => alu_res
                                      );

    set_status: process(alu_res) is
    begin
        if (alu_res = (others => '0')) then
            status(Z) <= '1';
        end if;
        status(S) <= alu_res(alu_res'high);
    end process set_status;

    alu_b <= b_reg when ctrl_alu_b = '0' else
             pc;

    alu_c <= c_reg when ctrl_alu_c = '0' else
             imm_reg;

    mdr_out <= b_reg;

end architecture rtl;
